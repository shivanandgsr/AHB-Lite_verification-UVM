class environment extends UVM_env;
`uvm_component_utils(environment)
  
  
